module MealyPattern(
	input        clock,
	input        i,
	output [1:0] o
);

// TODO Implementierung

endmodule

module MealyPatternTestbench();

	// TODO Input Stimuli

	MealyPattern machine(.clock(XXX), .i(XXX), .o(XXX));

	// TODO Überprüfe Ausgaben

endmodule

